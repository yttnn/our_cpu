typedef struct packed {
  logic lw;
  logic add;
  logic sub;
  logic addi;
} instructions;