module memory (

);
  
endmodule