typedef struct packed {
  logic lw;
  logic add;
} instructions;