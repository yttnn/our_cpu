typedef struct packed {
  logic lw;
  logic add;
  logic sub;
} instructions;